module axi_rw(
    
);