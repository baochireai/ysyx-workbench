module axi_rw(
    //pre_pc&&ifu
    //lsu&&wb
        
);