module ForwardUnit (
    input
);

endmodule