module top(
	input a,b,
	output f
);

assign f=a^b;

endmodule
